// Grant De La Campa
//
// mux4x1.v, 4x1 multiplexor, gate synthesis
//
// how to compile: ~changw/ivl/bin/iverilog mux2x1.v
// how to run: ./a.out

module MuxMod(s0, s1, d0, d1, d2, d3, o);
   input s0, s1, d0, d1, d2, d3;
   output o;

   wire s0_inv, s1_inv, and0, and_o, and1, and_1, and2, and_2, and3, and_3, or0, or1; // additional needed wires

   not(s0_inv, s0);
   not(s1_inv, s1);
   and(and0, s1_inv, s0_inv);
   and(and_0, and0, d0);
   and(and1, s1_inv, s0);
   and(and_1, and1, d1);
   and(and2, s1, s0_inv);
   and(and_2, and2, d2);
   and(and3, s1, s0);
   and(and_3, and3, d3);
   or(or0, and_0, and_1);
   or(or1, or0, and_2);
   or(o, or1, and_3);
   
endmodule

module TestMod;
   reg s0, s1, d0, d1, d2, d3;
   wire o;

   MuxMod my_mux(s0, s1, d0, d1, d2, d3, o);

//  initial #8 $finish; // end at $time 8

   initial begin
      $display("Time\ts0\ts1\td0\td1\td2\td3\to");
      $display("---------------------------------");
      $monitor("%0d\t%b\t%b\t%b\t%b\t%b\t%b\t%b", $time, s0, s1, d0, d1, d2, d3, o);
   end

   initial begin
      s0 = 0; s1 = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 0;   //000000
      #1;                      
      s0 = 0; s1 = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 1;   //000001
      #1; 
      s0 = 0; s1 = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 0;   //000010
      #1;                      
      s0 = 0; s1 = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 1;   //000011
      #1;                      
      s0 = 0; s1 = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 0;   //000100
      #1;                      
      s0 = 0; s1 = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 1;   //000101
      #1;                      
      s0 = 0; s1 = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 0;   //000110
      #1;                      
      s0 = 0; s1 = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 1;   //000111
      #1;                      
      s0 = 0; s1 = 0; d0 = 1; d1 = 0; d2 = 0; d3 = 0;   //001000
      #1;                      
      s0 = 0; s1 = 0; d0 = 1; d1 = 0; d2 = 0; d3 = 1;   //001001
      #1;                      
      s0 = 0; s1 = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 0;   //001010
      #1;                      
      s0 = 0; s1 = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 1;   //001011
      #1;                      
      s0 = 0; s1 = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 0;   //001100
      #1;                      
      s0 = 0; s1 = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 1;   //001101
      #1;
      s0 = 0; s1 = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 0;   //001110
      #1;       
      s0 = 0; s1 = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 1;   //001111
      #1;  
      s0 = 0; s1 = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 0;   //010000
      #1;                      
      s0 = 0; s1 = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 1;   //010001
      #1; 
      s0 = 0; s1 = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 0;   //010010
      #1;                      
      s0 = 0; s1 = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 1;   //010011
      #1;                      
      s0 = 0; s1 = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 0;   //010100
      #1;                      
      s0 = 0; s1 = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 1;   //010101
      #1;                    
      s0 = 0; s1 = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 0;   //010110
      #1;                      
      s0 = 0; s1 = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 1;   //010111
      #1;                      
      s0 = 0; s1 = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 0;   //011000
      #1;                      
      s0 = 0; s1 = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 1;   //011001
      #1;                      
      s0 = 0; s1 = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 0;   //011010
      #1;                      
      s0 = 0; s1 = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 1;   //011011
      #1;                      
      s0 = 0; s1 = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 0;   //011100
      #1;                      
      s0 = 0; s1 = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 1;   //011101
      #1;
      s0 = 0; s1 = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 0;   //011110
      #1;       
      s0 = 0; s1 = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 1;   //011111
      #1; 
      s0 = 1; s1 = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 0;   //100000
      #1;                      
      s0 = 1; s1 = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 1;   //100001
      #1; 
      s0 = 1; s1 = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 0;   //100010
      #1;                      
      s0 = 1; s1 = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 1;   //100011
      #1;                      
      s0 = 1; s1 = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 0;   //100100
      #1;                      
      s0 = 1; s1 = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 1;   //100101
      #1;                      
      s0 = 1; s1 = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 0;   //100110
      #1;                      
      s0 = 1; s1 = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 1;   //100111
      #1;                      
      s0 = 1; s1 = 0; d0 = 1; d1 = 0; d2 = 0; d3 = 0;   //101000
      #1;                      
      s0 = 1; s1 = 0; d0 = 1; d1 = 0; d2 = 0; d3 = 1;   //101001
      #1;                      
      s0 = 1; s1 = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 0;   //101010
      #1;                      
      s0 = 1; s1 = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 1;   //101011
      #1;                      
      s0 = 1; s1 = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 0;   //101100
      #1;                      
      s0 = 1; s1 = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 1;   //101101
      #1;
      s0 = 1; s1 = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 0;   //101110
      #1;       
      s0 = 1; s1 = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 1;   //101111
      #1;  
      s0 = 1; s1 = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 0;   //110000
      #1;                      
      s0 = 1; s1 = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 1;   //110001
      #1; 
      s0 = 1; s1 = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 0;   //110010
      #1;                      
      s0 = 1; s1 = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 1;   //110011
      #1;                      
      s0 = 1; s1 = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 0;   //110100
      #1;                      
      s0 = 1; s1 = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 1;   //110101
      #1;                    
      s0 = 1; s1 = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 0;   //110110
      #1;                      
      s0 = 1; s1 = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 1;   //110111
      #1;                      
      s0 = 1; s1 = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 0;   //111000
      #1;                      
      s0 = 1; s1 = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 1;   //111001
      #1;                      
      s0 = 1; s1 = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 0;   //111010
      #1;                      
      s0 = 1; s1 = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 1;   //111011
      #1;                      
      s0 = 1; s1 = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 0;   //111100
      #1;                      
      s0 = 1; s1 = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 1;   //111101
      #1;
      s0 = 1; s1 = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 0;   //111110
      #1;                            
      s0 = 1; s1 = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 1;   //111111
   end
endmodule